module top_module (
    input clk,
    input resetn,
    input [1:0] byteena,
    input [15:0] d,
    output reg [15:0] q
);
    wire [7:0] upper, lower;
    assign upper = d[15:8];
    assign lower = d[7:0];
    
    always @ (posedge clk) begin
        if (!resetn)
            q <= 16'b0;
        else begin
            if (byteena[0])
                q[7:0] <= d[7:0];
            if (byteena[1])
                q[15:8] <= d[15:8];
        end

    end

                
                

endmodule
